// The first verilog program to print "Hello World!"
module helloworld;
  initial begin;
    $display("Hello World!");
  end
endmodule
