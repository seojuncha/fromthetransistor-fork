module sram (
  input clk,
  input rst,
  input rd_en,   // read enable
  input wr_en,   // write enable
  input [15:0] address,
  input [31:0] data_in,
  output reg [31:0] data_out
);
  reg [31:0] memory [0:16383];

  // test fetch process only
  // explicitely copy a binary file into a current working directory.
  // initial begin
  //   $readmemb("little-mov.bin", memory);
  // end

  always @(posedge clk or negedge rst) begin
    if (!rst) begin
      memory <= 0;
      data_out <= 0;
    end else begin
      if (wr_en)
        memory[address] <= data_in;
      if (rd_en)
        data_out <= memory[address];
    end
  end

endmodule
