module bypass(
  input input_signal, 
  output output_signal
);
  assign output_signal = input_signal;
endmodule
