module not_child(
  input a,
  output not_a
);
  assign not_a = ~a;

endmodule
